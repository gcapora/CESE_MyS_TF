-- Archivo: cfa_seno.vhd
-- Autor:   Guillermo Caporaletti
-- Resumen: Conversor Fase-Amplitud para un NCO senoidal.
--          Trabajo Final del curso de CLP, CESE, FIUBA, Co18.
-- Fecha:   Junio 2023

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cfa_seno is
    generic (
        Q_BITS_DATO     : positive := 12;       -- Número de bits de cada dato-valor de salida (de 1 a 12)
        N_BITS_MUESTRAS : positive := 10        -- Bits necesario para las N muestras de señal por período
                                                -- 2^N_BITS_MUESTRAS debe ser >= 1024
    );
    port (
        reset_i  : in  std_logic;
        fase_i   : in  std_logic_vector(N_BITS_MUESTRAS - 1 downto 0);
        seno_o   : out std_logic_vector(Q_BITS_DATO - 1 downto 0)
    );
end entity cfa_seno;

architecture cfa_seno_arq of cfa_seno is
    constant Q_BITS_TDB : positive := 12;       -- Bits almacenados en la TdB
    constant N_MUESTRAS : positive := 1024;     -- Cantidad de muestras por período de señal 
    type tdb_type is array (0 to N_MUESTRAS - 1) of std_logic_vector(Q_BITS_TDB - 1 downto 0);
    constant tdb_seno   : tdb_type := (
        "011111111111", "100000001100", "100000011000", "100000100101", "100000110001", "100000111110", "100001001010", "100001010111", 
        "100001100011", "100001110000", "100001111101", "100010001001", "100010010110", "100010100010", "100010101111", "100010111011", 
        "100011001000", "100011010100", "100011100001", "100011101101", "100011111010", "100100000110", "100100010011", "100100011111", 
        "100100101011", "100100111000", "100101000100", "100101010001", "100101011101", "100101101001", "100101110110", "100110000010", 
        "100110001110", "100110011011", "100110100111", "100110110011", "100111000000", "100111001100", "100111011000", "100111100100", 
        "100111110001", "100111111101", "101000001001", "101000010101", "101000100001", "101000101101", "101000111001", "101001000101", 
        "101001010001", "101001011101", "101001101001", "101001110101", "101010000001", "101010001101", "101010011001", "101010100101", 
        "101010110001", "101010111101", "101011001000", "101011010100", "101011100000", "101011101100", "101011110111", "101100000011", 
        "101100001111", "101100011010", "101100100110", "101100110001", "101100111101", "101101001000", "101101010100", "101101011111", 
        "101101101010", "101101110110", "101110000001", "101110001100", "101110011000", "101110100011", "101110101110", "101110111001", 
        "101111000100", "101111001111", "101111011010", "101111100101", "101111110000", "101111111011", "110000000110", "110000010001", 
        "110000011100", "110000100110", "110000110001", "110000111100", "110001000110", "110001010001", "110001011100", "110001100110", 
        "110001110001", "110001111011", "110010000101", "110010010000", "110010011010", "110010100100", "110010101110", "110010111001", 
        "110011000011", "110011001101", "110011010111", "110011100001", "110011101011", "110011110101", "110011111110", "110100001000", 
        "110100010010", "110100011100", "110100100101", "110100101111", "110100111000", "110101000010", "110101001011", "110101010101", 
        "110101011110", "110101100111", "110101110001", "110101111010", "110110000011", "110110001100", "110110010101", "110110011110", 
        "110110100111", "110110110000", "110110111000", "110111000001", "110111001010", "110111010011", "110111011011", "110111100100", 
        "110111101100", "110111110101", "110111111101", "111000000101", "111000001101", "111000010110", "111000011110", "111000100110", 
        "111000101110", "111000110110", "111000111110", "111001000101", "111001001101", "111001010101", "111001011100", "111001100100", 
        "111001101100", "111001110011", "111001111010", "111010000010", "111010001001", "111010010000", "111010010111", "111010011110", 
        "111010100101", "111010101100", "111010110011", "111010111010", "111011000001", "111011001000", "111011001110", "111011010101", 
        "111011011011", "111011100010", "111011101000", "111011101110", "111011110101", "111011111011", "111100000001", "111100000111", 
        "111100001101", "111100010011", "111100011000", "111100011110", "111100100100", "111100101001", "111100101111", "111100110101", 
        "111100111010", "111100111111", "111101000101", "111101001010", "111101001111", "111101010100", "111101011001", "111101011110", 
        "111101100011", "111101100111", "111101101100", "111101110001", "111101110101", "111101111010", "111101111110", "111110000011", 
        "111110000111", "111110001011", "111110001111", "111110010011", "111110010111", "111110011011", "111110011111", "111110100011", 
        "111110100110", "111110101010", "111110101101", "111110110001", "111110110100", "111110111000", "111110111011", "111110111110", 
        "111111000001", "111111000100", "111111000111", "111111001010", "111111001101", "111111001111", "111111010010", "111111010101", 
        "111111010111", "111111011010", "111111011100", "111111011110", "111111100000", "111111100010", "111111100100", "111111100110", 
        "111111101000", "111111101010", "111111101100", "111111101110", "111111101111", "111111110001", "111111110010", "111111110011", 
        "111111110101", "111111110110", "111111110111", "111111111000", "111111111001", "111111111010", "111111111011", "111111111011", 
        "111111111100", "111111111101", "111111111101", "111111111110", "111111111110", "111111111110", "111111111110", "111111111110", 
        "111111111111", "111111111110", "111111111110", "111111111110", "111111111110", "111111111110", "111111111101", "111111111101", 
        "111111111100", "111111111011", "111111111011", "111111111010", "111111111001", "111111111000", "111111110111", "111111110110", 
        "111111110101", "111111110011", "111111110010", "111111110001", "111111101111", "111111101110", "111111101100", "111111101010", 
        "111111101000", "111111100110", "111111100100", "111111100010", "111111100000", "111111011110", "111111011100", "111111011010", 
        "111111010111", "111111010101", "111111010010", "111111001111", "111111001101", "111111001010", "111111000111", "111111000100", 
        "111111000001", "111110111110", "111110111011", "111110111000", "111110110100", "111110110001", "111110101101", "111110101010", 
        "111110100110", "111110100011", "111110011111", "111110011011", "111110010111", "111110010011", "111110001111", "111110001011", 
        "111110000111", "111110000011", "111101111110", "111101111010", "111101110101", "111101110001", "111101101100", "111101100111", 
        "111101100011", "111101011110", "111101011001", "111101010100", "111101001111", "111101001010", "111101000101", "111100111111", 
        "111100111010", "111100110101", "111100101111", "111100101001", "111100100100", "111100011110", "111100011000", "111100010011", 
        "111100001101", "111100000111", "111100000001", "111011111011", "111011110101", "111011101110", "111011101000", "111011100010", 
        "111011011011", "111011010101", "111011001110", "111011001000", "111011000001", "111010111010", "111010110011", "111010101100", 
        "111010100101", "111010011110", "111010010111", "111010010000", "111010001001", "111010000010", "111001111010", "111001110011", 
        "111001101100", "111001100100", "111001011100", "111001010101", "111001001101", "111001000101", "111000111110", "111000110110", 
        "111000101110", "111000100110", "111000011110", "111000010110", "111000001101", "111000000101", "110111111101", "110111110101", 
        "110111101100", "110111100100", "110111011011", "110111010011", "110111001010", "110111000001", "110110111000", "110110110000", 
        "110110100111", "110110011110", "110110010101", "110110001100", "110110000011", "110101111010", "110101110001", "110101100111", 
        "110101011110", "110101010101", "110101001011", "110101000010", "110100111000", "110100101111", "110100100101", "110100011100", 
        "110100010010", "110100001000", "110011111110", "110011110101", "110011101011", "110011100001", "110011010111", "110011001101", 
        "110011000011", "110010111001", "110010101110", "110010100100", "110010011010", "110010010000", "110010000101", "110001111011", 
        "110001110001", "110001100110", "110001011100", "110001010001", "110001000110", "110000111100", "110000110001", "110000100110", 
        "110000011100", "110000010001", "110000000110", "101111111011", "101111110000", "101111100101", "101111011010", "101111001111", 
        "101111000100", "101110111001", "101110101110", "101110100011", "101110011000", "101110001100", "101110000001", "101101110110", 
        "101101101010", "101101011111", "101101010100", "101101001000", "101100111101", "101100110001", "101100100110", "101100011010", 
        "101100001111", "101100000011", "101011110111", "101011101100", "101011100000", "101011010100", "101011001000", "101010111101", 
        "101010110001", "101010100101", "101010011001", "101010001101", "101010000001", "101001110101", "101001101001", "101001011101", 
        "101001010001", "101001000101", "101000111001", "101000101101", "101000100001", "101000010101", "101000001001", "100111111101", 
        "100111110001", "100111100100", "100111011000", "100111001100", "100111000000", "100110110011", "100110100111", "100110011011", 
        "100110001110", "100110000010", "100101110110", "100101101001", "100101011101", "100101010001", "100101000100", "100100111000", 
        "100100101011", "100100011111", "100100010011", "100100000110", "100011111010", "100011101101", "100011100001", "100011010100", 
        "100011001000", "100010111011", "100010101111", "100010100010", "100010010110", "100010001001", "100001111101", "100001110000", 
        "100001100011", "100001010111", "100001001010", "100000111110", "100000110001", "100000100101", "100000011000", "100000001100", 
        "011111111111", "011111110010", "011111100110", "011111011001", "011111001101", "011111000000", "011110110100", "011110100111", 
        "011110011011", "011110001110", "011110000001", "011101110101", "011101101000", "011101011100", "011101001111", "011101000011", 
        "011100110110", "011100101010", "011100011101", "011100010001", "011100000100", "011011111000", "011011101011", "011011011111", 
        "011011010011", "011011000110", "011010111010", "011010101101", "011010100001", "011010010101", "011010001000", "011001111100", 
        "011001110000", "011001100011", "011001010111", "011001001011", "011000111110", "011000110010", "011000100110", "011000011010", 
        "011000001101", "011000000001", "010111110101", "010111101001", "010111011101", "010111010001", "010111000101", "010110111001", 
        "010110101101", "010110100001", "010110010101", "010110001001", "010101111101", "010101110001", "010101100101", "010101011001", 
        "010101001101", "010101000001", "010100110110", "010100101010", "010100011110", "010100010010", "010100000111", "010011111011", 
        "010011101111", "010011100100", "010011011000", "010011001101", "010011000001", "010010110110", "010010101010", "010010011111", 
        "010010010100", "010010001000", "010001111101", "010001110010", "010001100110", "010001011011", "010001010000", "010001000101", 
        "010000111010", "010000101111", "010000100100", "010000011001", "010000001110", "010000000011", "001111111000", "001111101101", 
        "001111100010", "001111011000", "001111001101", "001111000010", "001110111000", "001110101101", "001110100010", "001110011000", 
        "001110001101", "001110000011", "001101111001", "001101101110", "001101100100", "001101011010", "001101010000", "001101000101", 
        "001100111011", "001100110001", "001100100111", "001100011101", "001100010011", "001100001001", "001100000000", "001011110110", 
        "001011101100", "001011100010", "001011011001", "001011001111", "001011000110", "001010111100", "001010110011", "001010101001", 
        "001010100000", "001010010111", "001010001101", "001010000100", "001001111011", "001001110010", "001001101001", "001001100000", 
        "001001010111", "001001001110", "001001000110", "001000111101", "001000110100", "001000101011", "001000100011", "001000011010", 
        "001000010010", "001000001001", "001000000001", "000111111001", "000111110001", "000111101000", "000111100000", "000111011000", 
        "000111010000", "000111001000", "000111000000", "000110111001", "000110110001", "000110101001", "000110100010", "000110011010", 
        "000110010010", "000110001011", "000110000100", "000101111100", "000101110101", "000101101110", "000101100111", "000101100000", 
        "000101011001", "000101010010", "000101001011", "000101000100", "000100111101", "000100110110", "000100110000", "000100101001", 
        "000100100011", "000100011100", "000100010110", "000100010000", "000100001001", "000100000011", "000011111101", "000011110111", 
        "000011110001", "000011101011", "000011100110", "000011100000", "000011011010", "000011010101", "000011001111", "000011001001", 
        "000011000100", "000010111111", "000010111001", "000010110100", "000010101111", "000010101010", "000010100101", "000010100000", 
        "000010011011", "000010010111", "000010010010", "000010001101", "000010001001", "000010000100", "000010000000", "000001111011", 
        "000001110111", "000001110011", "000001101111", "000001101011", "000001100111", "000001100011", "000001011111", "000001011011", 
        "000001011000", "000001010100", "000001010001", "000001001101", "000001001010", "000001000110", "000001000011", "000001000000", 
        "000000111101", "000000111010", "000000110111", "000000110100", "000000110001", "000000101111", "000000101100", "000000101001", 
        "000000100111", "000000100100", "000000100010", "000000100000", "000000011110", "000000011100", "000000011010", "000000011000", 
        "000000010110", "000000010100", "000000010010", "000000010000", "000000001111", "000000001101", "000000001100", "000000001011", 
        "000000001001", "000000001000", "000000000111", "000000000110", "000000000101", "000000000100", "000000000011", "000000000011", 
        "000000000010", "000000000001", "000000000001", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
        "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000001", "000000000001", 
        "000000000010", "000000000011", "000000000011", "000000000100", "000000000101", "000000000110", "000000000111", "000000001000", 
        "000000001001", "000000001011", "000000001100", "000000001101", "000000001111", "000000010000", "000000010010", "000000010100", 
        "000000010110", "000000011000", "000000011010", "000000011100", "000000011110", "000000100000", "000000100010", "000000100100", 
        "000000100111", "000000101001", "000000101100", "000000101111", "000000110001", "000000110100", "000000110111", "000000111010", 
        "000000111101", "000001000000", "000001000011", "000001000110", "000001001010", "000001001101", "000001010001", "000001010100", 
        "000001011000", "000001011011", "000001011111", "000001100011", "000001100111", "000001101011", "000001101111", "000001110011", 
        "000001110111", "000001111011", "000010000000", "000010000100", "000010001001", "000010001101", "000010010010", "000010010111", 
        "000010011011", "000010100000", "000010100101", "000010101010", "000010101111", "000010110100", "000010111001", "000010111111", 
        "000011000100", "000011001001", "000011001111", "000011010101", "000011011010", "000011100000", "000011100110", "000011101011", 
        "000011110001", "000011110111", "000011111101", "000100000011", "000100001001", "000100010000", "000100010110", "000100011100", 
        "000100100011", "000100101001", "000100110000", "000100110110", "000100111101", "000101000100", "000101001011", "000101010010", 
        "000101011001", "000101100000", "000101100111", "000101101110", "000101110101", "000101111100", "000110000100", "000110001011", 
        "000110010010", "000110011010", "000110100010", "000110101001", "000110110001", "000110111001", "000111000000", "000111001000", 
        "000111010000", "000111011000", "000111100000", "000111101000", "000111110001", "000111111001", "001000000001", "001000001001", 
        "001000010010", "001000011010", "001000100011", "001000101011", "001000110100", "001000111101", "001001000110", "001001001110", 
        "001001010111", "001001100000", "001001101001", "001001110010", "001001111011", "001010000100", "001010001101", "001010010111", 
        "001010100000", "001010101001", "001010110011", "001010111100", "001011000110", "001011001111", "001011011001", "001011100010", 
        "001011101100", "001011110110", "001100000000", "001100001001", "001100010011", "001100011101", "001100100111", "001100110001", 
        "001100111011", "001101000101", "001101010000", "001101011010", "001101100100", "001101101110", "001101111001", "001110000011", 
        "001110001101", "001110011000", "001110100010", "001110101101", "001110111000", "001111000010", "001111001101", "001111011000", 
        "001111100010", "001111101101", "001111111000", "010000000011", "010000001110", "010000011001", "010000100100", "010000101111", 
        "010000111010", "010001000101", "010001010000", "010001011011", "010001100110", "010001110010", "010001111101", "010010001000", 
        "010010010100", "010010011111", "010010101010", "010010110110", "010011000001", "010011001101", "010011011000", "010011100100", 
        "010011101111", "010011111011", "010100000111", "010100010010", "010100011110", "010100101010", "010100110110", "010101000001", 
        "010101001101", "010101011001", "010101100101", "010101110001", "010101111101", "010110001001", "010110010101", "010110100001", 
        "010110101101", "010110111001", "010111000101", "010111010001", "010111011101", "010111101001", "010111110101", "011000000001", 
        "011000001101", "011000011010", "011000100110", "011000110010", "011000111110", "011001001011", "011001010111", "011001100011", 
        "011001110000", "011001111100", "011010001000", "011010010101", "011010100001", "011010101101", "011010111010", "011011000110", 
        "011011010011", "011011011111", "011011101011", "011011111000", "011100000100", "011100010001", "011100011101", "011100101010", 
        "011100110110", "011101000011", "011101001111", "011101011100", "011101101000", "011101110101", "011110000001", "011110001110", 
        "011110011011", "011110100111", "011110110100", "011111000000", "011111001101", "011111011001", "011111100110", "011111110010" 
     );

    signal dato : std_logic_vector(Q_BITS_TDB - 1 downto 0);
    
begin

    process (fase_i, reset_i)
    begin
        if reset_i = '1' then
            dato <= (others => '0');
        else 
            dato <= tdb_seno(to_integer(unsigned(fase_i)));
        end if;
    end process;

    -- Puede ocurrir que se desee una salida con menos bots de cuantización.
    -- Por eso la diferencia entre Q_BITS_TDB y Q_BITS_DATO
    seno_o <= dato(Q_BITS_TDB-1 downto Q_BITS_TDB-Q_BITS_DATO);
    
end architecture cfa_seno_arq;
